/*
 * Calcula o CRC de data, compara com o crc recebido 
 * e coloca a resultado da compara��o em result
*/

module checksum (
	input  [7:0] data,	//Dado
	input  [7:0] crc,	//CRC
	output result		//Resultado
);

endmodule