// architecture.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module architecture (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n, // reset.reset_n
		output wire  uart_write,    //  uart.write
		input  wire  uart_read      //      .read
	);

	wire  [31:0] nios_data_master_readdata;                            // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                         // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                         // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [16:0] nios_data_master_address;                             // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                          // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                               // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                           // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                     // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                  // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [16:0] nios_instruction_master_address;                      // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                         // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire         mm_interconnect_0_arbitro_avalon_slave_0_chipselect;  // mm_interconnect_0:arbitro_avalon_slave_0_chipselect -> arbitro:chipselect
	wire  [31:0] mm_interconnect_0_arbitro_avalon_slave_0_readdata;    // arbitro:readdata -> mm_interconnect_0:arbitro_avalon_slave_0_readdata
	wire         mm_interconnect_0_arbitro_avalon_slave_0_read;        // mm_interconnect_0:arbitro_avalon_slave_0_read -> arbitro:read
	wire   [3:0] mm_interconnect_0_arbitro_avalon_slave_0_byteenable;  // mm_interconnect_0:arbitro_avalon_slave_0_byteenable -> arbitro:byteenable
	wire         mm_interconnect_0_arbitro_avalon_slave_0_write;       // mm_interconnect_0:arbitro_avalon_slave_0_write -> arbitro:write
	wire  [31:0] mm_interconnect_0_arbitro_avalon_slave_0_writedata;   // mm_interconnect_0:arbitro_avalon_slave_0_writedata -> arbitro:writedata
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;      // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;   // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;   // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;       // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;          // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;    // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;         // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;     // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;               // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                 // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [12:0] mm_interconnect_0_memory_s1_address;                  // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;               // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                    // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                    // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         irq_mapper_receiver0_irq;                             // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_irq_irq;                                         // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [arbitro:resetn, irq_mapper:reset, jtag:rst_n, memory:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [memory:reset_req, nios:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                       // nios:debug_reset_request -> rst_controller:reset_in1

	arbitro #(
		.uart_clock_bit (5208),
		.key            (9'b000110111)
	) arbitro (
		.resetn     (~rst_controller_reset_out_reset),                     //    clock_reset.reset_n
		.write      (mm_interconnect_0_arbitro_avalon_slave_0_write),      // avalon_slave_0.write
		.read       (mm_interconnect_0_arbitro_avalon_slave_0_read),       //               .read
		.chipselect (mm_interconnect_0_arbitro_avalon_slave_0_chipselect), //               .chipselect
		.byteenable (mm_interconnect_0_arbitro_avalon_slave_0_byteenable), //               .byteenable
		.writedata  (mm_interconnect_0_arbitro_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_arbitro_avalon_slave_0_readdata),   //               .readdata
		.clock      (clk_clk),                                             //     clock_sink.clk
		.tx         (uart_write),                                          //    conduit_end.write
		.rx         (uart_read)                                            //               .read
	);

	architecture_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	architecture_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	architecture_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	architecture_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                            (clk_clk),                                              //                          clk_clk.clk
		.nios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address               (nios_data_master_address),                             //                 nios_data_master.address
		.nios_data_master_waitrequest           (nios_data_master_waitrequest),                         //                                 .waitrequest
		.nios_data_master_byteenable            (nios_data_master_byteenable),                          //                                 .byteenable
		.nios_data_master_read                  (nios_data_master_read),                                //                                 .read
		.nios_data_master_readdata              (nios_data_master_readdata),                            //                                 .readdata
		.nios_data_master_write                 (nios_data_master_write),                               //                                 .write
		.nios_data_master_writedata             (nios_data_master_writedata),                           //                                 .writedata
		.nios_data_master_debugaccess           (nios_data_master_debugaccess),                         //                                 .debugaccess
		.nios_instruction_master_address        (nios_instruction_master_address),                      //          nios_instruction_master.address
		.nios_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                  //                                 .waitrequest
		.nios_instruction_master_read           (nios_instruction_master_read),                         //                                 .read
		.nios_instruction_master_readdata       (nios_instruction_master_readdata),                     //                                 .readdata
		.arbitro_avalon_slave_0_write           (mm_interconnect_0_arbitro_avalon_slave_0_write),       //           arbitro_avalon_slave_0.write
		.arbitro_avalon_slave_0_read            (mm_interconnect_0_arbitro_avalon_slave_0_read),        //                                 .read
		.arbitro_avalon_slave_0_readdata        (mm_interconnect_0_arbitro_avalon_slave_0_readdata),    //                                 .readdata
		.arbitro_avalon_slave_0_writedata       (mm_interconnect_0_arbitro_avalon_slave_0_writedata),   //                                 .writedata
		.arbitro_avalon_slave_0_byteenable      (mm_interconnect_0_arbitro_avalon_slave_0_byteenable),  //                                 .byteenable
		.arbitro_avalon_slave_0_chipselect      (mm_interconnect_0_arbitro_avalon_slave_0_chipselect),  //                                 .chipselect
		.jtag_avalon_jtag_slave_address         (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //           jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write           (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                 .write
		.jtag_avalon_jtag_slave_read            (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                 .read
		.jtag_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                 .readdata
		.jtag_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                 .writedata
		.jtag_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                 .waitrequest
		.jtag_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                 .chipselect
		.memory_s1_address                      (mm_interconnect_0_memory_s1_address),                  //                        memory_s1.address
		.memory_s1_write                        (mm_interconnect_0_memory_s1_write),                    //                                 .write
		.memory_s1_readdata                     (mm_interconnect_0_memory_s1_readdata),                 //                                 .readdata
		.memory_s1_writedata                    (mm_interconnect_0_memory_s1_writedata),                //                                 .writedata
		.memory_s1_byteenable                   (mm_interconnect_0_memory_s1_byteenable),               //                                 .byteenable
		.memory_s1_chipselect                   (mm_interconnect_0_memory_s1_chipselect),               //                                 .chipselect
		.memory_s1_clken                        (mm_interconnect_0_memory_s1_clken),                    //                                 .clken
		.nios_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),       //             nios_debug_mem_slave.address
		.nios_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),         //                                 .write
		.nios_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),          //                                 .read
		.nios_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),      //                                 .readdata
		.nios_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),     //                                 .writedata
		.nios_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),    //                                 .byteenable
		.nios_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest),   //                                 .waitrequest
		.nios_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess)    //                                 .debugaccess
	);

	architecture_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
