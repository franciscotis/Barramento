/*
 * Implementa a parte de emissor, do protocolo RS232
*/

module uart_tx (
	input  clock,
	input  reset,
	input  [7:0] data,	//Byte a ser enviado
	input  enable,		//Habilitado para iniciar envio

	output reg active,	//Habilitado durante o envio
	output reg done,	//Habilitado para envio conclu�do
	output reg tx		//Pino externo de sa�da do uart
);

endmodule