/*
 * Calcula o CRC de data, compara com o crc recebido 
 * e coloca a resultado da compara��o em result
*/

module checksum (
	input  [15:0] data,	//Dado e CRC recebidos
	output result		//Resultado
);

endmodule