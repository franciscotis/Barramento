
module architecture (
	clk_clk,
	reset_reset_n,
	uart_write,
	uart_read);	

	input		clk_clk;
	input		reset_reset_n;
	output		uart_write;
	input		uart_read;
endmodule
