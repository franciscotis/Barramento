/*
 * 
*/

module fsm (
	input clock,
	input reset,
	input data_rx,
	input active_tx,
	input done_tx,
	input result_crc,
	input  entry,			// Ser� utilizado para a mudan�a de estados
	output reg enable_tx,
	output reg [7:0] sensor

	//Entradas e sa�das do uart RS232
	input  rx,	//Pino externo de entrada
	output tx	//Pino externo de sa�da
);

//Declara��o do m�dulo emissor UART
wire [7:0] i_data_tx;	//N�mero do sensor
wire i_enable_tx;	//Habilita o envio do byte
wire o_active_tx;	//Habilitado enquanto o byte est� sendo enviado
wire o_done_tx;		//Habilitado quando o byte foi enviado

//Declara��o do m�dulodo receptor UART
wire [15:0] o_data_rx;	//2 bytes recebidos
wire o_done_rx;		//Habilitado quando os 2 bytes s�o recebidos

//Declara��o do m�dulo de verica��o do CRC
wire o_result_crc;	//Resultado da verfica��o




parameter [2:0] A = 3'b000, //Nomes dos estados 
		B = 3'b001,
		C = 3'b010,
		D = 3'b011,
		E = 3'b100,
		F = 3'b101,
		G = 3'b111;

reg [1:0] state,next;

localparam 	STATE_1 = 3'b000, //Par�metros locais utilizados para a compara��o com a entrada
		STATE_2 = 3'b001,
		STATE_3 = 3'b010,
		STATE_4 = 3'b011,
		STATE_5 = 3'b100,
		STATE_6 = 3'b101,
		STATE_7 = 3'b111;

always @(posedge clock or negedge reset)
	if (!reset) state <= A;
	else 	    state <= next;


always @(state) begin
	next = 3'bx;
	result = 8'b00000000;

case(state)
	A: 
	if(entry == STATE_1) next = A;
	else if(entry == STATE_2) next = B;
	else if(entry == STATE_3) next = C;
	else if(entry == STATE_4) next = D;
	else if(entry == STATE_5) next = E;
	else if(entry == STATE_6) next = F;
	B:
	if(entry == STATE_1) next = A;
	else 
		uart_tx UART_TX (.clock(clock), .reset(~reset), .data(i_data_tx), .enable(i_enable_tx), 
		.active(o_active_tx), .done(o_done_tx), .tx(tx));
		#10;
		uart_rx UART_RX (.clock(clock), .reset(~reset), .rx(rx), .data(o_data_rx), .done(o_done_rx));	
		#5;
		checksum CHECKSUM (.data(o_data_rx[7:0]), .crc(o_data_rx[15:8]), .result(o_result_crc));
		assign result = o_result_crc;
	C:
	if(entry == STATE_1) next = A;
	else 
		uart_tx UART_TX (.clock(clock), .reset(~reset), .data(i_data_tx), .enable(i_enable_tx), 
		.active(o_active_tx), .done(o_done_tx), .tx(tx));
		#10;
		uart_rx UART_RX (.clock(clock), .reset(~reset), .rx(rx), .data(o_data_rx), .done(o_done_rx));	
		#5;
		checksum CHECKSUM (.data(o_data_rx[7:0]), .crc(o_data_rx[15:8]), .result(o_result_crc));
		assign result = o_result_crc;
	D:
	if(entry == STATE_1) next = A;
	else 
		uart_tx UART_TX (.clock(clock), .reset(~reset), .data(i_data_tx), .enable(i_enable_tx), 
		.active(o_active_tx), .done(o_done_tx), .tx(tx));
		#10;
		uart_rx UART_RX (.clock(clock), .reset(~reset), .rx(rx), .data(o_data_rx), .done(o_done_rx));	
		#5;
		checksum CHECKSUM (.data(o_data_rx[7:0]), .crc(o_data_rx[15:8]), .result(o_result_crc));
		assign result = o_result_crc;
		
	E:
	if(entry == STATE_1) next = A;
	else 
		uart_tx UART_TX (.clock(clock), .reset(~reset), .data(i_data_tx), .enable(i_enable_tx), 
		.active(o_active_tx), .done(o_done_tx), .tx(tx));
		#10;
		uart_rx UART_RX (.clock(clock), .reset(~reset), .rx(rx), .data(o_data_rx), .done(o_done_rx));	
		#5;
		checksum CHECKSUM (.data(o_data_rx[7:0]), .crc(o_data_rx[15:8]), .result(o_result_crc));
		assign result = o_result_crc;
	F:
	if(entry == STATE_1) next = A;
	else 
		uart_tx UART_TX (.clock(clock), .reset(~reset), .data(i_data_tx), .enable(i_enable_tx), 
		.active(o_active_tx), .done(o_done_tx), .tx(tx));
		#10;
		uart_rx UART_RX (.clock(clock), .reset(~reset), .rx(rx), .data(o_data_rx), .done(o_done_rx));	
		#5;
		checksum CHECKSUM (.data(o_data_rx[7:0]), .crc(o_data_rx[15:8]), .result(o_result_crc));
		assign result = o_result_crc;

endcase
end


endmodule	